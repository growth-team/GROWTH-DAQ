library ieee, work;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package TestWaveform is

  type   Vector12Bits is array (natural range<>) of std_logic_vector(11 downto 0);
  constant TestWaveformGaus : Vector12Bits(599 downto 0) := (
        77 => conv_std_logic_vector(0, 12),
        78 => conv_std_logic_vector(1, 12),
        79 => conv_std_logic_vector(1, 12),
        80 => conv_std_logic_vector(1, 12),
        81 => conv_std_logic_vector(1, 12),
        82 => conv_std_logic_vector(1, 12),
        83 => conv_std_logic_vector(1, 12),
        84 => conv_std_logic_vector(1, 12),
        85 => conv_std_logic_vector(2, 12),
        86 => conv_std_logic_vector(2, 12),
        87 => conv_std_logic_vector(2, 12),
        88 => conv_std_logic_vector(2, 12),
        89 => conv_std_logic_vector(2, 12),
        90 => conv_std_logic_vector(3, 12),
        91 => conv_std_logic_vector(3, 12),
        92 => conv_std_logic_vector(3, 12),
        93 => conv_std_logic_vector(4, 12),
        94 => conv_std_logic_vector(4, 12),
        95 => conv_std_logic_vector(4, 12),
        96 => conv_std_logic_vector(5, 12),
        97 => conv_std_logic_vector(5, 12),
        98 => conv_std_logic_vector(6, 12),
        99 => conv_std_logic_vector(6, 12),
        100 => conv_std_logic_vector(7, 12),
        101 => conv_std_logic_vector(7, 12),
        102 => conv_std_logic_vector(8, 12),
        103 => conv_std_logic_vector(9, 12),
        104 => conv_std_logic_vector(10, 12),
        105 => conv_std_logic_vector(10, 12),
        106 => conv_std_logic_vector(11, 12),
        107 => conv_std_logic_vector(12, 12),
        108 => conv_std_logic_vector(13, 12),
        109 => conv_std_logic_vector(14, 12),
        110 => conv_std_logic_vector(15, 12),
        111 => conv_std_logic_vector(16, 12),
        112 => conv_std_logic_vector(18, 12),
        113 => conv_std_logic_vector(19, 12),
        114 => conv_std_logic_vector(20, 12),
        115 => conv_std_logic_vector(22, 12),
        116 => conv_std_logic_vector(23, 12),
        117 => conv_std_logic_vector(25, 12),
        118 => conv_std_logic_vector(27, 12),
        119 => conv_std_logic_vector(28, 12),
        120 => conv_std_logic_vector(30, 12),
        121 => conv_std_logic_vector(32, 12),
        122 => conv_std_logic_vector(35, 12),
        123 => conv_std_logic_vector(37, 12),
        124 => conv_std_logic_vector(39, 12),
        125 => conv_std_logic_vector(42, 12),
        126 => conv_std_logic_vector(44, 12),
        127 => conv_std_logic_vector(47, 12),
        128 => conv_std_logic_vector(50, 12),
        129 => conv_std_logic_vector(53, 12),
        130 => conv_std_logic_vector(56, 12),
        131 => conv_std_logic_vector(59, 12),
        132 => conv_std_logic_vector(62, 12),
        133 => conv_std_logic_vector(66, 12),
        134 => conv_std_logic_vector(70, 12),
        135 => conv_std_logic_vector(73, 12),
        136 => conv_std_logic_vector(77, 12),
        137 => conv_std_logic_vector(81, 12),
        138 => conv_std_logic_vector(85, 12),
        139 => conv_std_logic_vector(90, 12),
        140 => conv_std_logic_vector(94, 12),
        141 => conv_std_logic_vector(99, 12),
        142 => conv_std_logic_vector(104, 12),
        143 => conv_std_logic_vector(109, 12),
        144 => conv_std_logic_vector(114, 12),
        145 => conv_std_logic_vector(119, 12),
        146 => conv_std_logic_vector(124, 12),
        147 => conv_std_logic_vector(130, 12),
        148 => conv_std_logic_vector(135, 12),
        149 => conv_std_logic_vector(141, 12),
        150 => conv_std_logic_vector(147, 12),
        151 => conv_std_logic_vector(153, 12),
        152 => conv_std_logic_vector(159, 12),
        153 => conv_std_logic_vector(165, 12),
        154 => conv_std_logic_vector(171, 12),
        155 => conv_std_logic_vector(177, 12),
        156 => conv_std_logic_vector(184, 12),
        157 => conv_std_logic_vector(190, 12),
        158 => conv_std_logic_vector(197, 12),
        159 => conv_std_logic_vector(204, 12),
        160 => conv_std_logic_vector(210, 12),
        161 => conv_std_logic_vector(217, 12),
        162 => conv_std_logic_vector(224, 12),
        163 => conv_std_logic_vector(231, 12),
        164 => conv_std_logic_vector(238, 12),
        165 => conv_std_logic_vector(245, 12),
        166 => conv_std_logic_vector(251, 12),
        167 => conv_std_logic_vector(258, 12),
        168 => conv_std_logic_vector(265, 12),
        169 => conv_std_logic_vector(272, 12),
        170 => conv_std_logic_vector(279, 12),
        171 => conv_std_logic_vector(285, 12),
        172 => conv_std_logic_vector(292, 12),
        173 => conv_std_logic_vector(298, 12),
        174 => conv_std_logic_vector(305, 12),
        175 => conv_std_logic_vector(311, 12),
        176 => conv_std_logic_vector(317, 12),
        177 => conv_std_logic_vector(323, 12),
        178 => conv_std_logic_vector(329, 12),
        179 => conv_std_logic_vector(335, 12),
        180 => conv_std_logic_vector(340, 12),
        181 => conv_std_logic_vector(346, 12),
        182 => conv_std_logic_vector(351, 12),
        183 => conv_std_logic_vector(356, 12),
        184 => conv_std_logic_vector(361, 12),
        185 => conv_std_logic_vector(365, 12),
        186 => conv_std_logic_vector(369, 12),
        187 => conv_std_logic_vector(373, 12),
        188 => conv_std_logic_vector(377, 12),
        189 => conv_std_logic_vector(381, 12),
        190 => conv_std_logic_vector(384, 12),
        191 => conv_std_logic_vector(387, 12),
        192 => conv_std_logic_vector(389, 12),
        193 => conv_std_logic_vector(392, 12),
        194 => conv_std_logic_vector(394, 12),
        195 => conv_std_logic_vector(396, 12),
        196 => conv_std_logic_vector(397, 12),
        197 => conv_std_logic_vector(398, 12),
        198 => conv_std_logic_vector(399, 12),
        199 => conv_std_logic_vector(399, 12),
        200 => conv_std_logic_vector(400, 12),
        201 => conv_std_logic_vector(399, 12),
        202 => conv_std_logic_vector(399, 12),
        203 => conv_std_logic_vector(398, 12),
        204 => conv_std_logic_vector(397, 12),
        205 => conv_std_logic_vector(396, 12),
        206 => conv_std_logic_vector(394, 12),
        207 => conv_std_logic_vector(392, 12),
        208 => conv_std_logic_vector(389, 12),
        209 => conv_std_logic_vector(387, 12),
        210 => conv_std_logic_vector(384, 12),
        211 => conv_std_logic_vector(381, 12),
        212 => conv_std_logic_vector(377, 12),
        213 => conv_std_logic_vector(373, 12),
        214 => conv_std_logic_vector(369, 12),
        215 => conv_std_logic_vector(365, 12),
        216 => conv_std_logic_vector(361, 12),
        217 => conv_std_logic_vector(356, 12),
        218 => conv_std_logic_vector(351, 12),
        219 => conv_std_logic_vector(346, 12),
        220 => conv_std_logic_vector(340, 12),
        221 => conv_std_logic_vector(335, 12),
        222 => conv_std_logic_vector(329, 12),
        223 => conv_std_logic_vector(323, 12),
        224 => conv_std_logic_vector(317, 12),
        225 => conv_std_logic_vector(311, 12),
        226 => conv_std_logic_vector(305, 12),
        227 => conv_std_logic_vector(298, 12),
        228 => conv_std_logic_vector(292, 12),
        229 => conv_std_logic_vector(285, 12),
        230 => conv_std_logic_vector(279, 12),
        231 => conv_std_logic_vector(272, 12),
        232 => conv_std_logic_vector(265, 12),
        233 => conv_std_logic_vector(258, 12),
        234 => conv_std_logic_vector(251, 12),
        235 => conv_std_logic_vector(245, 12),
        236 => conv_std_logic_vector(238, 12),
        237 => conv_std_logic_vector(231, 12),
        238 => conv_std_logic_vector(224, 12),
        239 => conv_std_logic_vector(217, 12),
        240 => conv_std_logic_vector(210, 12),
        241 => conv_std_logic_vector(204, 12),
        242 => conv_std_logic_vector(197, 12),
        243 => conv_std_logic_vector(190, 12),
        244 => conv_std_logic_vector(184, 12),
        245 => conv_std_logic_vector(177, 12),
        246 => conv_std_logic_vector(171, 12),
        247 => conv_std_logic_vector(165, 12),
        248 => conv_std_logic_vector(159, 12),
        249 => conv_std_logic_vector(153, 12),
        250 => conv_std_logic_vector(147, 12),
        251 => conv_std_logic_vector(141, 12),
        252 => conv_std_logic_vector(135, 12),
        253 => conv_std_logic_vector(130, 12),
        254 => conv_std_logic_vector(124, 12),
        255 => conv_std_logic_vector(119, 12),
        256 => conv_std_logic_vector(114, 12),
        257 => conv_std_logic_vector(109, 12),
        258 => conv_std_logic_vector(104, 12),
        259 => conv_std_logic_vector(99, 12),
        260 => conv_std_logic_vector(94, 12),
        261 => conv_std_logic_vector(90, 12),
        262 => conv_std_logic_vector(85, 12),
        263 => conv_std_logic_vector(81, 12),
        264 => conv_std_logic_vector(77, 12),
        265 => conv_std_logic_vector(73, 12),
        266 => conv_std_logic_vector(70, 12),
        267 => conv_std_logic_vector(66, 12),
        268 => conv_std_logic_vector(62, 12),
        269 => conv_std_logic_vector(59, 12),
        270 => conv_std_logic_vector(56, 12),
        271 => conv_std_logic_vector(53, 12),
        272 => conv_std_logic_vector(50, 12),
        273 => conv_std_logic_vector(47, 12),
        274 => conv_std_logic_vector(44, 12),
        275 => conv_std_logic_vector(42, 12),
        276 => conv_std_logic_vector(39, 12),
        277 => conv_std_logic_vector(37, 12),
        278 => conv_std_logic_vector(35, 12),
        279 => conv_std_logic_vector(32, 12),
        280 => conv_std_logic_vector(30, 12),
        281 => conv_std_logic_vector(28, 12),
        282 => conv_std_logic_vector(27, 12),
        283 => conv_std_logic_vector(25, 12),
        284 => conv_std_logic_vector(23, 12),
        285 => conv_std_logic_vector(22, 12),
        286 => conv_std_logic_vector(20, 12),
        287 => conv_std_logic_vector(19, 12),
        288 => conv_std_logic_vector(18, 12),
        289 => conv_std_logic_vector(16, 12),
        290 => conv_std_logic_vector(15, 12),
        291 => conv_std_logic_vector(14, 12),
        292 => conv_std_logic_vector(13, 12),
        293 => conv_std_logic_vector(12, 12),
        294 => conv_std_logic_vector(11, 12),
        295 => conv_std_logic_vector(10, 12),
        296 => conv_std_logic_vector(10, 12),
        297 => conv_std_logic_vector(9, 12),
        298 => conv_std_logic_vector(8, 12),
        299 => conv_std_logic_vector(7, 12),
        300 => conv_std_logic_vector(7, 12),
        301 => conv_std_logic_vector(6, 12),
        302 => conv_std_logic_vector(6, 12),
        303 => conv_std_logic_vector(5, 12),
        304 => conv_std_logic_vector(5, 12),
        305 => conv_std_logic_vector(4, 12),
        306 => conv_std_logic_vector(4, 12),
        307 => conv_std_logic_vector(4, 12),
        308 => conv_std_logic_vector(3, 12),
        309 => conv_std_logic_vector(3, 12),
        310 => conv_std_logic_vector(3, 12),
        311 => conv_std_logic_vector(2, 12),
        312 => conv_std_logic_vector(2, 12),
        313 => conv_std_logic_vector(2, 12),
        314 => conv_std_logic_vector(2, 12),
        315 => conv_std_logic_vector(2, 12),
        316 => conv_std_logic_vector(1, 12),
        317 => conv_std_logic_vector(1, 12),
        318 => conv_std_logic_vector(1, 12),
        319 => conv_std_logic_vector(1, 12),
        320 => conv_std_logic_vector(1, 12),
        321 => conv_std_logic_vector(1, 12),
        322 => conv_std_logic_vector(1, 12),
        323 => conv_std_logic_vector(0, 12),
        others =>  (others => '0')
  );

end TestWaveform;
